`include "constants.v"

module 