//(c) Chris Adams 2015 - Uinversity of Leeds.

//Constants

`define OSC_DEPTH 16
`define OSC_AMP_MAX 65536

//NUmber of words in the half sine memory
`define HALF_SINE_WORDS 65536