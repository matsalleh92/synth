//(c) Chris Adams 2015 - Uinversity of Leeds.

//Top level for my really bad synth

module synth (input clk);
	//OTB oscillator_tb;
	
	oscillator_tb OTB();
endmodule